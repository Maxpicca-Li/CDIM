module d_cache #(
    parameter LEN_LINE = 6,  // 64 Bytes
    parameter LEN_INDEX = 6, // 64 lines
    parameter NR_WAYS = 2,
    parameter SIZE_STORE_BUFFER = 8
) (
    input               clk,
    input               rst,
    // to cpu
    input               stallM,
    output              dstall,
    input        [31:0] E_mem_pa, // only used for match bram
    input        [31:0] M_mem_pa,
    input        [31:0] M_fence_addr, // used for fence
    input               M_fence_d, // fence address reuse the M_memva. Note: we shouldn't raise M_fence_en with M_mem_en.
    input               M_mem_en,
    input               M_mem_write,
    input               M_mem_uncached,
    input        [ 3:0] M_wmask,
    input         [1:0] M_mem_size,
    input        [31:0] M_wdata,
    output       [31:0] M_rdata,
    // to axi
    output logic [31:0] araddr,
    output logic [ 7:0] arlen,
    output logic [ 2:0] arsize,
    output logic        arvalid,
    input               arready,
    input  [31:0]       rdata,
    input               rlast,
    input               rvalid,
    output logic        rready,
    output logic [31:0] awaddr,
    output logic  [7:0] awlen,
    output logic  [2:0] awsize,
    output logic        awvalid,
    input               awready,
    output logic [31:0] wdata,
    output logic [3: 0] wstrb,
    output logic        wlast,
    output logic        wvalid,
    input               wready,
    input               bvalid,
    output              bready
);

// defines

localparam LEN_PER_WAY = LEN_LINE + LEN_INDEX;
localparam LEN_TAG = 32 - LEN_LINE - LEN_INDEX;
localparam LEN_BRAM_ADDR = LEN_LINE - 3 + LEN_INDEX;
localparam NR_LINES = 1 << LEN_INDEX;
localparam NR_WORDS = 1 << (LEN_LINE - 2);

typedef struct packed {
    logic [LEN_TAG-1:0] tag;
} dcache_tag;

typedef struct packed {
    logic [NR_WAYS-1:0] valid;
    logic [NR_WAYS-1:0] dirty;
    logic LRU;
    // Note: If NR_WAYS > 2, we should implement pseudo-LRU or LFSR.
} dcache_meta;

enum { IDLE, UNCACHED_READ, CACHE_WRITEBACK, CACHE_REPLACE, SAVE_RESULT } dcache_status;

// metadata
dcache_meta meta [NR_LINES-1:0];

// mmio store buffer
typedef struct packed {
    logic [31:0]    waddr;
    logic [1:0]     wsize;
    logic [3:0]     wstrb;
    logic [31:0]    wdata; // note: data should place at correct place. (like axi)
} store_buffer_entry;

typedef struct packed {
    logic [$clog2(SIZE_STORE_BUFFER)-1:0] ptr_begin;
    logic [$clog2(SIZE_STORE_BUFFER)-1:0] ptr_end;
    logic axi_busy;
} store_buffer_control;

store_buffer_entry store_buffer[SIZE_STORE_BUFFER-1:0];
store_buffer_control store_buffer_ctrl;
logic current_mmio_write_saved;
wire store_buffer_has_next = store_buffer_ctrl.ptr_begin != store_buffer_ctrl.ptr_end;
wire store_buffer_busy = store_buffer_has_next | store_buffer_ctrl.axi_busy;
wire store_buffer_full = (store_buffer_ctrl.ptr_end + 3'd1) == store_buffer_ctrl.ptr_begin;

// replace & fence control
wire [LEN_PER_WAY-1:LEN_LINE]   fence_line_addr = M_fence_addr[LEN_PER_WAY-1:LEN_LINE];
logic [LEN_LINE-1:2] axi_rcnt; // cache -> axi_w cnt
logic [LEN_LINE-1:2] axi_wcnt; // axi_r -> cache cnt
logic [LEN_PER_WAY-1:2] bram_replace_addr;
logic [LEN_PER_WAY-1:2] bram_read_ready_addr;
logic [LEN_PER_WAY-1:2] bram_replace_write_addr;
logic [$clog2(NR_WORDS):0] bram_replace_cnt; // cnt itself can be send to axi (by mux cache_data[i] and bram_r_buffer), cnt - 1 can be read from bram_r_buffer
logic [31:0] bram_r_buffer [NR_WORDS-1:0];
logic bram_use_replace_addr;
logic bram_data_valid;
logic fence_working;
logic aw_handshake;
logic replace_writeback;
wire fence_way = meta[fence_line_addr].dirty[1] ? 1'b1 : 1'b0;
// TODO: If we changed NR_WAYS, we should add judge to each way

logic tag_wea[NR_WAYS-1:0];
logic [3:0] bram_replace_wea [NR_WAYS-1:0];

wire [3:0] data_wea [NR_WAYS-1:0]; // assign at generate

dcache_tag tag_ram_wdata;

// dcache bram
wire [31:LEN_PER_WAY] addr_tag = M_mem_pa[31:LEN_PER_WAY];
wire bram_addr_choose = dstall | stallM; // 1: M_mem_pa or M_fence_addr, 0: E_mem_pa

// FIXME: fix M_fence_addr
wire [LEN_PER_WAY-1:2]          bram_word_addr = bram_use_replace_addr ? bram_replace_addr : (bram_addr_choose ? M_mem_pa[LEN_PER_WAY-1:2] : E_mem_pa[LEN_PER_WAY-1:2]);
wire [LEN_PER_WAY-1:LEN_LINE]   bram_line_addr = bram_use_replace_addr ? bram_replace_addr[LEN_PER_WAY-1:LEN_LINE] : (bram_addr_choose ? M_mem_pa[LEN_PER_WAY-1:LEN_LINE] : E_mem_pa[LEN_PER_WAY-1:LEN_LINE]);

wire [LEN_PER_WAY-1:2] tag_read_addr = bram_word_addr;
wire [LEN_PER_WAY-1:2] data_read_addr = bram_word_addr;
wire [LEN_PER_WAY-1:2] data_write_addr = bram_use_replace_addr ? bram_replace_write_addr : M_mem_pa[LEN_PER_WAY-1:2];

wire data_bram_wdata_sel = dcache_status == CACHE_REPLACE; // 1: axi rdata, 0: M_wdata
wire [31:0] data_bram_wdata = data_bram_wdata_sel ? rdata : M_wdata;

wire [31:0] cache_data [NR_WAYS-1:0];
dcache_tag cache_tag[NR_WAYS-1:0];

wire [NR_WAYS-1:0] tag_compare_valid;
wire cache_hit = |tag_compare_valid;

wire cache_hit_available = cache_hit && !M_mem_uncached;

// stall control
wire mmio_read_stall = M_mem_en && M_mem_uncached && !M_mem_write && dcache_status != SAVE_RESULT;
wire mmio_write_stall = (M_mem_en && M_mem_uncached && M_mem_write && (dcache_status != IDLE || store_buffer_full) );
wire cached_stall = M_mem_en & (!M_mem_uncached) & !cache_hit;
wire fence_stall = M_fence_d && dcache_status != SAVE_RESULT;

// Note: If NR_WAYS > 2, we should mux one hot from tag_compare_valid;
wire d_cache_sel = tag_compare_valid[1];

wire [LEN_PER_WAY-1:LEN_LINE] pa_line_addr = M_mem_pa[LEN_PER_WAY-1:LEN_LINE];

assign dstall = dcache_status == IDLE ? ((cached_stall | mmio_read_stall | mmio_write_stall) | M_fence_d) : (dcache_status != SAVE_RESULT);

logic [31:0] saved_rdata;

// forward last stored data in data bram
logic [LEN_PER_WAY-1:2] last_line_addr; // two way shared
logic [31:0] last_wea [NR_WAYS-1:0]; // assume only write one way at a time
logic [31:0] last_wdata; // two way shared
wire [31:0] cache_data_forward [NR_WAYS-1:0];

assign M_rdata = dcache_status == SAVE_RESULT ? saved_rdata : cache_data_forward[d_cache_sel];

// generate bram
genvar i;
generate
    for (i=0;i<NR_WAYS;i++) begin
        dual_port_bram_bw8 #(.LEN_DATA(32),.LEN_ADDR(LEN_PER_WAY-2)) d_data
        (
            .clka   (clk),
            .clkb   (clk),
            .ena    (1'b1),
            .enb    (1'b1),
            .addra  (data_write_addr),
            .dina   (data_bram_wdata),
            .wea    (data_wea[i]),
            .addrb  (bram_word_addr),
            .doutb  (cache_data[i])
        );
        dual_port_bram_nobw #(.LEN_DATA(LEN_TAG),.LEN_ADDR(LEN_PER_WAY-LEN_LINE)) d_tag
        (
            .clka   (clk),
            .clkb   (clk),
            .ena    (1'b1),
            .enb    (1'b1),
            .addra  (bram_replace_addr[LEN_PER_WAY-1:LEN_LINE]),
            .dina   (tag_ram_wdata),
            .wea    (tag_wea[i]),
            .addrb  (bram_line_addr),
            .doutb  (cache_tag[i])
        );
        assign tag_compare_valid[i] = cache_tag[i].tag == addr_tag && meta[pa_line_addr].valid[i];
        assign cache_data_forward[i] = (last_wea[i] & last_wdata) | (cache_data[i] & (~last_wea[i]));
        assign data_wea[i] = (tag_compare_valid[i] && M_mem_en && M_mem_write && !M_mem_uncached && dcache_status == IDLE) ? M_wmask :  bram_replace_wea[i];
        always_ff @(posedge clk) begin
            if (rst) begin
                last_wea[i] <= 0;
            end
            else begin
                last_wea[i] <= {{8{data_wea[i][3]}},{8{data_wea[i][2]}},{8{data_wea[i][1]}},{8{data_wea[i][0]}}};
            end
        end
    end
endgenerate
// save last_line_addr
always_ff @(posedge clk) begin
    if (rst) begin
        last_line_addr <= 0;
        last_wdata <= 0;
    end
    else begin
        last_line_addr <= bram_word_addr;
        last_wdata <= data_bram_wdata;
    end
end

// axi bready
assign bready = 1'b1;


always_ff @(posedge clk) begin
    if (rst) begin
        // clear store buffer
        store_buffer_ctrl <= 0;
        current_mmio_write_saved <= 0;
        // clear replace ctrl
        axi_rcnt <= 0;
        axi_wcnt <= 0;
        bram_replace_addr <= 0;
        bram_read_ready_addr <= 0;
        bram_replace_cnt <= 0;
        bram_r_buffer <= '{default: '0};
        bram_use_replace_addr <= 0;
        bram_replace_write_addr <= 0;
        bram_data_valid <= 0;
        fence_working <= 0;
        aw_handshake <= 0;
        replace_writeback <= 0;
        tag_wea <= '{default: '0};
        bram_replace_wea <= '{default: '0};
        tag_ram_wdata <= 0;
        // clear saved rdata
        saved_rdata <= 0;
        // clear axi
        araddr <= 0;
        arlen <= 0;
        arsize <= 0;
        arvalid <= 0;
        rready <= 0;
        awaddr <= 0;
        awlen <= 0;
        awsize <= 0;
        awvalid <= 0;
        wdata <= 0;
        wstrb <= 0;
        wlast <= 0;
        wvalid <= 0;
    end
    else begin
        // store buffer
        if (store_buffer_busy) begin
            if (store_buffer_ctrl.axi_busy) begin // To implement SC memory ordering, if store buffer busy, axi is unseable.
                if (awvalid & awready) begin
                    awvalid <= 0;
                end
                if (wvalid & wready) begin
                    if (store_buffer_has_next) begin
                        awaddr <= store_buffer[store_buffer_ctrl.ptr_begin].waddr;
                        awlen <= 0;
                        awsize <= {1'd0,store_buffer[store_buffer_ctrl.ptr_begin].wsize};
                        awvalid <= 1'b1;
                        wdata <= store_buffer[store_buffer_ctrl.ptr_begin].wdata;
                        wstrb <= store_buffer[store_buffer_ctrl.ptr_begin].wstrb;
                        wlast <= 1'b1;
                        wvalid <= 1'b1;
                        store_buffer_ctrl.ptr_begin <= store_buffer_ctrl.ptr_begin + 3'd1;
                    end
                    else begin
                        wvalid <= 0;
                        wlast <= 0;
                        store_buffer_ctrl.axi_busy <= 1'b0;
                    end
                end
            end
            else begin
                awaddr <= store_buffer[store_buffer_ctrl.ptr_begin].waddr;
                awlen <= 0;
                awsize <= {1'd0,store_buffer[store_buffer_ctrl.ptr_begin].wsize};
                awvalid <= 1'b1;
                wdata <= store_buffer[store_buffer_ctrl.ptr_begin].wdata;
                wstrb <= store_buffer[store_buffer_ctrl.ptr_begin].wstrb;
                wlast <= 1'b1;
                wvalid <= 1'b1;
                store_buffer_ctrl.ptr_begin <= store_buffer_ctrl.ptr_begin + 3'd1;
                store_buffer_ctrl.axi_busy <= 1'b1;
            end
        end
        case (dcache_status)
            IDLE: begin
                if (M_mem_en) begin
                    if (M_mem_uncached) begin
                        if (M_mem_write) begin
                            if (!store_buffer_full && !current_mmio_write_saved) begin
                                store_buffer[store_buffer_ctrl.ptr_end] <= '{
                                    waddr: M_mem_pa,
                                    wsize: M_mem_size,
                                    wstrb: M_wmask,
                                    wdata: M_wdata
                                };
                                store_buffer_ctrl.ptr_end <= store_buffer_ctrl.ptr_end + 3'd1;
                                current_mmio_write_saved <= 1'b1;
                            end
                            if (!dstall && !stallM) begin
                                current_mmio_write_saved <= 1'b0;
                            end
                        end
                        else begin // mmio read
                            if (!store_buffer_busy) begin
                                araddr <= M_mem_pa;
                                arlen <= 0;
                                arsize <= {1'b0, M_mem_size};
                                arvalid <= 1'b1;
                                dcache_status <= UNCACHED_READ;
                                rready <= 1'b1;
                            end // if store buffer busy, read will stop at IDLE but stall pipeline.
                        end
                    end
                    else begin
                        if (!cache_hit) begin

                        end
                        else begin
                            if (!dstall && !stallM) begin
                                // Update LRU
                                meta[pa_line_addr].LRU <= ~d_cache_sel;
                            end
                        end
                    end
                end
                else if (M_fence_d) begin
                    if (|meta[fence_line_addr].dirty) begin
                        dcache_status <= CACHE_WRITEBACK;
                        axi_rcnt <= 0;
                        axi_wcnt <= 0;
                        bram_replace_addr <= {M_fence_addr[LEN_PER_WAY-1:LEN_LINE],{LEN_LINE-2{1'b0}}};
                        bram_read_ready_addr <= {M_fence_addr[LEN_PER_WAY-1:LEN_LINE],{LEN_LINE-2{1'b0}}};
                        bram_replace_cnt <= 0;
                        bram_use_replace_addr <= 1'b1;
                        bram_data_valid <= 0;
                    end
                    else if (|meta[fence_line_addr].valid) begin
                        meta[fence_line_addr].valid <= 0;
                        dcache_status <= SAVE_RESULT;
                    end
                end
            end
            UNCACHED_READ: begin
                if (arvalid && arready) begin
                    arvalid <= 1'b0;
                end
                if (rvalid) begin
                    saved_rdata <= rdata;
                    dcache_status <= SAVE_RESULT;
                end
            end
            CACHE_WRITEBACK: begin // CACHE Instruction
                if (fence_working) begin
                    if (bram_replace_addr[LEN_LINE-1:2] != NR_WORDS - 1) begin
                        bram_replace_addr <= bram_replace_addr + 1;
                    end
                    bram_read_ready_addr <= bram_replace_addr;
                    bram_r_buffer[bram_read_ready_addr[LEN_LINE-1:2]] <= cache_data[fence_way];
                    if (!aw_handshake) begin
                        awaddr <= {cache_tag[fence_way].tag,fence_line_addr,{LEN_LINE{1'b0}}};
                        awlen <= NR_WORDS - 1;
                        awsize <= 3'd2;
                        awvalid <= 1'b1;
                        wdata <= cache_data[fence_way];
                        wstrb <= 4'b1111;
                        wlast <= NR_WORDS == 1 ? 1'b1 : 1'b0;
                        wvalid <= 1'b1;
                        aw_handshake <= 1'b1;
                    end
                    if (awvalid & awready) begin
                        awvalid <= 1'b0;
                    end
                    if (wvalid & wready) begin
                        if (wlast) begin
                            wvalid <= 1'b0;
                            meta[fence_line_addr].dirty[fence_way] <= 1'b0;
                            fence_working <= 1'b0;
                            bram_use_replace_addr <= 1'b0;
                            dcache_status <= IDLE;
                        end
                        else begin
                            wdata <= ((axi_wcnt + 1'b1) == bram_read_ready_addr[LEN_LINE-1:2]) ? cache_data[fence_way] : bram_r_buffer[axi_wcnt + 1'b1];
                            axi_wcnt <= axi_wcnt + 1;
                            if ({1'b0,axi_wcnt} + 1'b1 == NR_WORDS - 1) begin
                                wlast <= 1'b1;
                            end
                        end
                    end
                end
                else begin
                    aw_handshake <= 1'b0;
                    fence_working <= 1'b1;
                    bram_replace_addr[LEN_LINE-1:2] <= bram_replace_addr[LEN_LINE-1:2] + 1;
                    // transfer [addr + 1], and receive [addr].
                end
            end
            CACHE_REPLACE: begin
                
            end
            SAVE_RESULT: begin
                if (!dstall && !stallM) begin
                    dcache_status <= IDLE;
                end
            end
        endcase
    end
end

endmodule
